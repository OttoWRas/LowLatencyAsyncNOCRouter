LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.math_real.ALL;
USE work.internals.ALL;
USE work.defs.ALL;

ENTITY router_top_tb IS
END ENTITY;

ARCHITECTURE impl OF router_top_tb IS
    DUT : router_top PORT MAP(
        ports
    );
BEGIN
END ARCHITECTURE;

